/* 

David Fritz and Brian Gordon 

VGA module, framebuffer, and signal generator

Memory map:

0xf0400000 - control register
0xf0400004 - frame buffer pointer

*/

module mod_vga(rst, clk, ie, de, iaddr, daddr, drw, din, iout, dout, rgb, hs, vs);
        input rst;
        input clk;
        input ie,de;
        input [31:0] iaddr, daddr;
        input drw;
        input [31:0] din;
        output [31:0] iout, dout;
        output [7:0] rgb;
	output hs, vs;

        /* by spec, the iout and dout signals must go hiZ when we're not using them */
        wire [31:0] idata, ddata;
        assign iout = ie ? idata : 32'hzzzzzzzz;
        assign dout = de ? ddata : 32'hzzzzzzzz;

        assign idata = 32'h00000000;

	wire [7:0] eff_rgb;
	wire [10:0] hcount, vcount;
	wire blank, fb_write;

	reg enable;
	reg [31:0] fb_pointer;
	
	/* the vga controller */
	vga_controller vga(clk, rst, hs, vs, blank, hcount, vcount);
	vga_sram_bypass bypass(clk, fb_pointer, hcount, vcount, eff_rgb);

	always @(negedge clk) begin
		if (drw && de) begin
			if (daddr == 32'h00000000)
				enable <= din[0];
			else if (daddr == 32'h00000004)
				fb_pointer <= din;
		end
	end			

	assign rgb = (blank) ? 0 : 
		     (enable) ? eff_rgb : 0;
endmodule

module vga_controller (clk, rst, hs, vs, blank, hcount, vcount);

  input             clk, rst;
  output 	        hs, vs;
  output reg 		  blank;
  output reg [10:0] hcount, vcount;
  reg        [10:0] hcounter, vcounter;
  
  parameter H_FRONTPORCH = 16;
  parameter H_BACKPORCH  = 48;
  parameter H_PULSEWIDTH = 96;
  parameter H_PERIOD     = 800;
  
  parameter V_FRONTPORCH = 10;
  parameter V_BACKPORCH  = 29;
  parameter V_PULSEWIDTH = 2;
  parameter V_PERIOD     = 521;
    
  assign hs = (hcounter < H_PULSEWIDTH) ? 0 : 1;
  assign vs = (vcounter < V_PULSEWIDTH) ? 0 : 1;
   
  always @(negedge clk) begin
	if (rst) begin
		hcount   = 0;
		vcount   = 0;
		hcounter = 0;
		vcounter = 0;
		blank    = 1;
	end
  
    // blank signal
    blank = (hcounter >= H_PULSEWIDTH + H_BACKPORCH && 
             hcounter <  H_PERIOD - H_FRONTPORCH &&
             vcounter >= V_PULSEWIDTH + V_BACKPORCH &&
             vcounter <  V_PERIOD - V_FRONTPORCH)
             ? 0 : 1;
             
    //hcount = (blank) ? 0 : hcount + 1;
    //Vcount = (blank) ? 0 : Vcount + 1;
             
    hcounter = hcounter + 1;
    if (hcounter == H_PERIOD) begin
      hcounter = 0;
      vcounter = (vcounter == V_PERIOD) ? 0 : vcounter + 1;
    end

    hcount = ((hcounter >= H_PULSEWIDTH + H_BACKPORCH) && 
              (hcounter <  H_PERIOD - H_FRONTPORCH))
              ? (hcounter - H_PULSEWIDTH) - H_BACKPORCH : 0;
              
    vcount = ((vcounter >= V_PULSEWIDTH + V_BACKPORCH) &&
              (vcounter <  V_PERIOD - V_FRONTPORCH))
              ? (vcounter - V_PULSEWIDTH) - V_BACKPORCH : 0;
    
  end
endmodule

module vga_sram_bypass (clk, fb_addr, hcount, vcount, rgb);
	input clk;
	input [31:0] fb_addr;
	input [10:0] hcount, vcount;
	output [7:0] rgb;

	reg [7:0] buffer [639:0]; /* our buffer */
	
	/* we use hcount to index into the buffer */
	assign rgb = buffer[hcount];

initial begin
buffer[0] = 0;
buffer[1] = 1;
buffer[2] = 2;
buffer[3] = 3;
buffer[4] = 4;
buffer[5] = 5;
buffer[6] = 6;
buffer[7] = 7;
buffer[8] = 8;
buffer[9] = 9;
buffer[10] = 10;
buffer[11] = 11;
buffer[12] = 12;
buffer[13] = 13;
buffer[14] = 14;
buffer[15] = 15;
buffer[16] = 16;
buffer[17] = 17;
buffer[18] = 18;
buffer[19] = 19;
buffer[20] = 20;
buffer[21] = 21;
buffer[22] = 22;
buffer[23] = 23;
buffer[24] = 24;
buffer[25] = 25;
buffer[26] = 26;
buffer[27] = 27;
buffer[28] = 28;
buffer[29] = 29;
buffer[30] = 30;
buffer[31] = 31;
buffer[32] = 32;
buffer[33] = 33;
buffer[34] = 34;
buffer[35] = 35;
buffer[36] = 36;
buffer[37] = 37;
buffer[38] = 38;
buffer[39] = 39;
buffer[40] = 40;
buffer[41] = 41;
buffer[42] = 42;
buffer[43] = 43;
buffer[44] = 44;
buffer[45] = 45;
buffer[46] = 46;
buffer[47] = 47;
buffer[48] = 48;
buffer[49] = 49;
buffer[50] = 50;
buffer[51] = 51;
buffer[52] = 52;
buffer[53] = 53;
buffer[54] = 54;
buffer[55] = 55;
buffer[56] = 56;
buffer[57] = 57;
buffer[58] = 58;
buffer[59] = 59;
buffer[60] = 60;
buffer[61] = 61;
buffer[62] = 62;
buffer[63] = 63;
buffer[64] = 64;
buffer[65] = 65;
buffer[66] = 66;
buffer[67] = 67;
buffer[68] = 68;
buffer[69] = 69;
buffer[70] = 70;
buffer[71] = 71;
buffer[72] = 72;
buffer[73] = 73;
buffer[74] = 74;
buffer[75] = 75;
buffer[76] = 76;
buffer[77] = 77;
buffer[78] = 78;
buffer[79] = 79;
buffer[80] = 80;
buffer[81] = 81;
buffer[82] = 82;
buffer[83] = 83;
buffer[84] = 84;
buffer[85] = 85;
buffer[86] = 86;
buffer[87] = 87;
buffer[88] = 88;
buffer[89] = 89;
buffer[90] = 90;
buffer[91] = 91;
buffer[92] = 92;
buffer[93] = 93;
buffer[94] = 94;
buffer[95] = 95;
buffer[96] = 96;
buffer[97] = 97;
buffer[98] = 98;
buffer[99] = 99;
buffer[100] = 100;
buffer[101] = 101;
buffer[102] = 102;
buffer[103] = 103;
buffer[104] = 104;
buffer[105] = 105;
buffer[106] = 106;
buffer[107] = 107;
buffer[108] = 108;
buffer[109] = 109;
buffer[110] = 110;
buffer[111] = 111;
buffer[112] = 112;
buffer[113] = 113;
buffer[114] = 114;
buffer[115] = 115;
buffer[116] = 116;
buffer[117] = 117;
buffer[118] = 118;
buffer[119] = 119;
buffer[120] = 120;
buffer[121] = 121;
buffer[122] = 122;
buffer[123] = 123;
buffer[124] = 124;
buffer[125] = 125;
buffer[126] = 126;
buffer[127] = 127;
buffer[128] = 128;
buffer[129] = 129;
buffer[130] = 130;
buffer[131] = 131;
buffer[132] = 132;
buffer[133] = 133;
buffer[134] = 134;
buffer[135] = 135;
buffer[136] = 136;
buffer[137] = 137;
buffer[138] = 138;
buffer[139] = 139;
buffer[140] = 140;
buffer[141] = 141;
buffer[142] = 142;
buffer[143] = 143;
buffer[144] = 144;
buffer[145] = 145;
buffer[146] = 146;
buffer[147] = 147;
buffer[148] = 148;
buffer[149] = 149;
buffer[150] = 150;
buffer[151] = 151;
buffer[152] = 152;
buffer[153] = 153;
buffer[154] = 154;
buffer[155] = 155;
buffer[156] = 156;
buffer[157] = 157;
buffer[158] = 158;
buffer[159] = 159;
buffer[160] = 160;
buffer[161] = 161;
buffer[162] = 162;
buffer[163] = 163;
buffer[164] = 164;
buffer[165] = 165;
buffer[166] = 166;
buffer[167] = 167;
buffer[168] = 168;
buffer[169] = 169;
buffer[170] = 170;
buffer[171] = 171;
buffer[172] = 172;
buffer[173] = 173;
buffer[174] = 174;
buffer[175] = 175;
buffer[176] = 176;
buffer[177] = 177;
buffer[178] = 178;
buffer[179] = 179;
buffer[180] = 180;
buffer[181] = 181;
buffer[182] = 182;
buffer[183] = 183;
buffer[184] = 184;
buffer[185] = 185;
buffer[186] = 186;
buffer[187] = 187;
buffer[188] = 188;
buffer[189] = 189;
buffer[190] = 190;
buffer[191] = 191;
buffer[192] = 192;
buffer[193] = 193;
buffer[194] = 194;
buffer[195] = 195;
buffer[196] = 196;
buffer[197] = 197;
buffer[198] = 198;
buffer[199] = 199;
buffer[200] = 200;
buffer[201] = 201;
buffer[202] = 202;
buffer[203] = 203;
buffer[204] = 204;
buffer[205] = 205;
buffer[206] = 206;
buffer[207] = 207;
buffer[208] = 208;
buffer[209] = 209;
buffer[210] = 210;
buffer[211] = 211;
buffer[212] = 212;
buffer[213] = 213;
buffer[214] = 214;
buffer[215] = 215;
buffer[216] = 216;
buffer[217] = 217;
buffer[218] = 218;
buffer[219] = 219;
buffer[220] = 220;
buffer[221] = 221;
buffer[222] = 222;
buffer[223] = 223;
buffer[224] = 224;
buffer[225] = 225;
buffer[226] = 226;
buffer[227] = 227;
buffer[228] = 228;
buffer[229] = 229;
buffer[230] = 230;
buffer[231] = 231;
buffer[232] = 232;
buffer[233] = 233;
buffer[234] = 234;
buffer[235] = 235;
buffer[236] = 236;
buffer[237] = 237;
buffer[238] = 238;
buffer[239] = 239;
buffer[240] = 240;
buffer[241] = 241;
buffer[242] = 242;
buffer[243] = 243;
buffer[244] = 244;
buffer[245] = 245;
buffer[246] = 246;
buffer[247] = 247;
buffer[248] = 248;
buffer[249] = 249;
buffer[250] = 250;
buffer[251] = 251;
buffer[252] = 252;
buffer[253] = 253;
buffer[254] = 254;
buffer[255] = 255;
buffer[256] = 0;
buffer[257] = 1;
buffer[258] = 2;
buffer[259] = 3;
buffer[260] = 4;
buffer[261] = 5;
buffer[262] = 6;
buffer[263] = 7;
buffer[264] = 8;
buffer[265] = 9;
buffer[266] = 10;
buffer[267] = 11;
buffer[268] = 12;
buffer[269] = 13;
buffer[270] = 14;
buffer[271] = 15;
buffer[272] = 16;
buffer[273] = 17;
buffer[274] = 18;
buffer[275] = 19;
buffer[276] = 20;
buffer[277] = 21;
buffer[278] = 22;
buffer[279] = 23;
buffer[280] = 24;
buffer[281] = 25;
buffer[282] = 26;
buffer[283] = 27;
buffer[284] = 28;
buffer[285] = 29;
buffer[286] = 30;
buffer[287] = 31;
buffer[288] = 32;
buffer[289] = 33;
buffer[290] = 34;
buffer[291] = 35;
buffer[292] = 36;
buffer[293] = 37;
buffer[294] = 38;
buffer[295] = 39;
buffer[296] = 40;
buffer[297] = 41;
buffer[298] = 42;
buffer[299] = 43;
buffer[300] = 44;
buffer[301] = 45;
buffer[302] = 46;
buffer[303] = 47;
buffer[304] = 48;
buffer[305] = 49;
buffer[306] = 50;
buffer[307] = 51;
buffer[308] = 52;
buffer[309] = 53;
buffer[310] = 54;
buffer[311] = 55;
buffer[312] = 56;
buffer[313] = 57;
buffer[314] = 58;
buffer[315] = 59;
buffer[316] = 60;
buffer[317] = 61;
buffer[318] = 62;
buffer[319] = 63;
buffer[320] = 64;
buffer[321] = 65;
buffer[322] = 66;
buffer[323] = 67;
buffer[324] = 68;
buffer[325] = 69;
buffer[326] = 70;
buffer[327] = 71;
buffer[328] = 72;
buffer[329] = 73;
buffer[330] = 74;
buffer[331] = 75;
buffer[332] = 76;
buffer[333] = 77;
buffer[334] = 78;
buffer[335] = 79;
buffer[336] = 80;
buffer[337] = 81;
buffer[338] = 82;
buffer[339] = 83;
buffer[340] = 84;
buffer[341] = 85;
buffer[342] = 86;
buffer[343] = 87;
buffer[344] = 88;
buffer[345] = 89;
buffer[346] = 90;
buffer[347] = 91;
buffer[348] = 92;
buffer[349] = 93;
buffer[350] = 94;
buffer[351] = 95;
buffer[352] = 96;
buffer[353] = 97;
buffer[354] = 98;
buffer[355] = 99;
buffer[356] = 100;
buffer[357] = 101;
buffer[358] = 102;
buffer[359] = 103;
buffer[360] = 104;
buffer[361] = 105;
buffer[362] = 106;
buffer[363] = 107;
buffer[364] = 108;
buffer[365] = 109;
buffer[366] = 110;
buffer[367] = 111;
buffer[368] = 112;
buffer[369] = 113;
buffer[370] = 114;
buffer[371] = 115;
buffer[372] = 116;
buffer[373] = 117;
buffer[374] = 118;
buffer[375] = 119;
buffer[376] = 120;
buffer[377] = 121;
buffer[378] = 122;
buffer[379] = 123;
buffer[380] = 124;
buffer[381] = 125;
buffer[382] = 126;
buffer[383] = 127;
buffer[384] = 128;
buffer[385] = 129;
buffer[386] = 130;
buffer[387] = 131;
buffer[388] = 132;
buffer[389] = 133;
buffer[390] = 134;
buffer[391] = 135;
buffer[392] = 136;
buffer[393] = 137;
buffer[394] = 138;
buffer[395] = 139;
buffer[396] = 140;
buffer[397] = 141;
buffer[398] = 142;
buffer[399] = 143;
buffer[400] = 144;
buffer[401] = 145;
buffer[402] = 146;
buffer[403] = 147;
buffer[404] = 148;
buffer[405] = 149;
buffer[406] = 150;
buffer[407] = 151;
buffer[408] = 152;
buffer[409] = 153;
buffer[410] = 154;
buffer[411] = 155;
buffer[412] = 156;
buffer[413] = 157;
buffer[414] = 158;
buffer[415] = 159;
buffer[416] = 160;
buffer[417] = 161;
buffer[418] = 162;
buffer[419] = 163;
buffer[420] = 164;
buffer[421] = 165;
buffer[422] = 166;
buffer[423] = 167;
buffer[424] = 168;
buffer[425] = 169;
buffer[426] = 170;
buffer[427] = 171;
buffer[428] = 172;
buffer[429] = 173;
buffer[430] = 174;
buffer[431] = 175;
buffer[432] = 176;
buffer[433] = 177;
buffer[434] = 178;
buffer[435] = 179;
buffer[436] = 180;
buffer[437] = 181;
buffer[438] = 182;
buffer[439] = 183;
buffer[440] = 184;
buffer[441] = 185;
buffer[442] = 186;
buffer[443] = 187;
buffer[444] = 188;
buffer[445] = 189;
buffer[446] = 190;
buffer[447] = 191;
buffer[448] = 192;
buffer[449] = 193;
buffer[450] = 194;
buffer[451] = 195;
buffer[452] = 196;
buffer[453] = 197;
buffer[454] = 198;
buffer[455] = 199;
buffer[456] = 200;
buffer[457] = 201;
buffer[458] = 202;
buffer[459] = 203;
buffer[460] = 204;
buffer[461] = 205;
buffer[462] = 206;
buffer[463] = 207;
buffer[464] = 208;
buffer[465] = 209;
buffer[466] = 210;
buffer[467] = 211;
buffer[468] = 212;
buffer[469] = 213;
buffer[470] = 214;
buffer[471] = 215;
buffer[472] = 216;
buffer[473] = 217;
buffer[474] = 218;
buffer[475] = 219;
buffer[476] = 220;
buffer[477] = 221;
buffer[478] = 222;
buffer[479] = 223;
buffer[480] = 224;
buffer[481] = 225;
buffer[482] = 226;
buffer[483] = 227;
buffer[484] = 228;
buffer[485] = 229;
buffer[486] = 230;
buffer[487] = 231;
buffer[488] = 232;
buffer[489] = 233;
buffer[490] = 234;
buffer[491] = 235;
buffer[492] = 236;
buffer[493] = 237;
buffer[494] = 238;
buffer[495] = 239;
buffer[496] = 240;
buffer[497] = 241;
buffer[498] = 242;
buffer[499] = 243;
buffer[500] = 244;
buffer[501] = 245;
buffer[502] = 246;
buffer[503] = 247;
buffer[504] = 248;
buffer[505] = 249;
buffer[506] = 250;
buffer[507] = 251;
buffer[508] = 252;
buffer[509] = 253;
buffer[510] = 254;
buffer[511] = 255;
buffer[512] = 0;
buffer[513] = 1;
buffer[514] = 2;
buffer[515] = 3;
buffer[516] = 4;
buffer[517] = 5;
buffer[518] = 6;
buffer[519] = 7;
buffer[520] = 8;
buffer[521] = 9;
buffer[522] = 10;
buffer[523] = 11;
buffer[524] = 12;
buffer[525] = 13;
buffer[526] = 14;
buffer[527] = 15;
buffer[528] = 16;
buffer[529] = 17;
buffer[530] = 18;
buffer[531] = 19;
buffer[532] = 20;
buffer[533] = 21;
buffer[534] = 22;
buffer[535] = 23;
buffer[536] = 24;
buffer[537] = 25;
buffer[538] = 26;
buffer[539] = 27;
buffer[540] = 28;
buffer[541] = 29;
buffer[542] = 30;
buffer[543] = 31;
buffer[544] = 32;
buffer[545] = 33;
buffer[546] = 34;
buffer[547] = 35;
buffer[548] = 36;
buffer[549] = 37;
buffer[550] = 38;
buffer[551] = 39;
buffer[552] = 40;
buffer[553] = 41;
buffer[554] = 42;
buffer[555] = 43;
buffer[556] = 44;
buffer[557] = 45;
buffer[558] = 46;
buffer[559] = 47;
buffer[560] = 48;
buffer[561] = 49;
buffer[562] = 50;
buffer[563] = 51;
buffer[564] = 52;
buffer[565] = 53;
buffer[566] = 54;
buffer[567] = 55;
buffer[568] = 56;
buffer[569] = 57;
buffer[570] = 58;
buffer[571] = 59;
buffer[572] = 60;
buffer[573] = 61;
buffer[574] = 62;
buffer[575] = 63;
buffer[576] = 64;
buffer[577] = 65;
buffer[578] = 66;
buffer[579] = 67;
buffer[580] = 68;
buffer[581] = 69;
buffer[582] = 70;
buffer[583] = 71;
buffer[584] = 72;
buffer[585] = 73;
buffer[586] = 74;
buffer[587] = 75;
buffer[588] = 76;
buffer[589] = 77;
buffer[590] = 78;
buffer[591] = 79;
buffer[592] = 80;
buffer[593] = 81;
buffer[594] = 82;
buffer[595] = 83;
buffer[596] = 84;
buffer[597] = 85;
buffer[598] = 86;
buffer[599] = 87;
buffer[600] = 88;
buffer[601] = 89;
buffer[602] = 90;
buffer[603] = 91;
buffer[604] = 92;
buffer[605] = 93;
buffer[606] = 94;
buffer[607] = 95;
buffer[608] = 96;
buffer[609] = 97;
buffer[610] = 98;
buffer[611] = 99;
buffer[612] = 100;
buffer[613] = 101;
buffer[614] = 102;
buffer[615] = 103;
buffer[616] = 104;
buffer[617] = 105;
buffer[618] = 106;
buffer[619] = 107;
buffer[620] = 108;
buffer[621] = 109;
buffer[622] = 110;
buffer[623] = 111;
buffer[624] = 112;
buffer[625] = 113;
buffer[626] = 114;
buffer[627] = 115;
buffer[628] = 116;
buffer[629] = 117;
buffer[630] = 118;
buffer[631] = 119;
buffer[632] = 120;
buffer[633] = 121;
buffer[634] = 122;
buffer[635] = 123;
buffer[636] = 124;
buffer[637] = 125;
buffer[638] = 126;
buffer[639] = 127;
end
endmodule

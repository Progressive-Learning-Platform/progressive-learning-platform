module bar;

 initial $display("lib/bar.v %l");

endmodule

module foo;

 initial $display("foo/foo.v %l");

endmodule

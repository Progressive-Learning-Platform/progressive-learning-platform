module foo1;

 initial $display("foo/foo1.v %l");

endmodule

module foo2;

 initial $display("foo/foo2.v %l");

endmodule

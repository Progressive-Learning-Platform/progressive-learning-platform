module xx;
 initial $display("hello world.");
endmodule

module adder;

 initial $display("lib/adder.v adder %l");

endmodule

module adder2;

 initial $display("lib/adder.v adder2 %l");

endmodule
